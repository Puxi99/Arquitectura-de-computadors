library ieee;
use ieee.std_logic_1164.all;

entity CPU is
    Port(
        clock,reset: in std_logic;
    )
end entity;

architecture behavior of CPU is
    begin
        
    end behavior;